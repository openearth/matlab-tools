netcdf netCDF4_tutorial_grid_lat_lon_curvilinear {
dimensions:
	col = 3 ;
	row = 5 ;
	time = 1 ;
	bounds = 4 ;
variables:
	double time(time) ;
		time:standard_name = "time" ;
		time:long_name = "time" ;
		time:units = "seconds since 1970-01-01 00-00-00" ;
		time:axis = "T" ;
	double lon(row, col) ;
		lon:_FillValue = 1.#QNAN000000000 ;
		lon:standard_name = "longitude" ;
		lon:long_name = "Longitude" ;
		lon:units = "degrees_east" ;
		lon:axis = "X" ;
		lon:grid_mapping = "projection" ;
		lon:actual_range = 2., 6. ;
		lon:bounds = "lon_bnds" ;
	double lat(row, col) ;
		lat:_FillValue = 1.#QNAN000000000 ;
		lat:standard_name = "latitude" ;
		lat:long_name = "Latitude" ;
		lat:units = "degrees_north" ;
		lat:axis = "Y" ;
		lat:grid_mapping = "projection" ;
		lat:actual_range = 50., 54. ;
		lat:bounds = "lat_bnds" ;
	int projection ;
		projection:name = "WGS 84" ;
		projection:epsg = 4326. ;
		projection:grid_mapping_name = "latitude_longitude" ;
		projection:semi_major_axis = 6378137. ;
		projection:semi_minor_axis = 6356752.31424783 ;
		projection:inverse_flattening = 298.2572236 ;
		projection:proj4_params = "+proj=longlat +ellps=WGS84 +datum=WGS84 +no_defs" ;
		projection:projection_name = "Latitude Longitude" ;
		projection:EPSG_code = "EPSG:4326" ;
	double lon_bnds(row, col, bounds) ;
		lon_bnds:_FillValue = 1.#QNAN000000000 ;
		lon_bnds:standard_name = "longitude" ;
		lon_bnds:long_name = "Longitude bounds" ;
		lon_bnds:units = "degrees_east" ;
		lon_bnds:actual_range = 1., 7. ;
	double lat_bnds(row, col, bounds) ;
		lat_bnds:_FillValue = 1.#QNAN000000000 ;
		lat_bnds:standard_name = "latitude" ;
		lat_bnds:long_name = "Latitude bounds" ;
		lat_bnds:units = "degrees_north" ;
		lat_bnds:actual_range = 49.5, 54.5 ;
	float depth(time, row, col) ;
		depth:_FillValue = 1.#QNAN0f ;
		depth:standard_name = "sea_floor_depth_below_geoid" ;
		depth:long_name = "bottom depth" ;
		depth:units = "m" ;
		depth:positive = "up" ;
		depth:actual_range = 1., 114. ;
		depth:grid_mapping = "projection" ;
		depth:coordinates = "lat lon" ;

// global attributes:
		:title = "ncwritetutorial_grid_lat_lon_curvilinear" ;
		:institution = "Deltares" ;
		:source = "X" ;
		:history = "$HeadURL: https://svn.oss.deltares.nl/repos/openearthtools/trunk/python/OpenEarthTools/openearthtools/io/netcdf/netCDF4_tutorial_grid_lat_lon_curvilinear.cdl $ $Id: netCDF4_tutorial_grid_lat_lon_curvilinear.cdl 8907 2013-07-10 12:39:16Z boer_g $" ;
		:references = "http://svn.oss.deltares.nl" ;
		:email = "X" ;
		:featureType = "Grid" ;
		:comment = "X" ;
		:version = "beta" ;
		:Conventions = "CF-1.6" ;
		:terms_for_use = "These data can be used freely for research purposes provided that the following source is acknowledged: Deltares" ;
		:disclaimer = "This data is made available in the hope that it will be useful, but WITHOUT ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE." ;
data:

 time = 946681200 ;

 lon =
  2, 4, 6,
  2, 4, 6,
  2, 4, 1.#QNAN,
  2, 4, 6,
  2, 4, 6 ;

 lat =
  50, 50, 50,
  51, 51, 51,
  52, 52, 1.#QNAN,
  53, 53, 53,
  54, 54, 54 ;

 projection = _ ;

 lon_bnds =
  1, 3, 3, 1,
  3, 5, 5, 3,
  5, 7, 7, 5,
  1, 3, 3, 1,
  3, 5, 5, 3,
  5, 7, 7, 5,
  1, 3, 3, 1,
  3, 5, 5, 3,
  5, 7, 7, 5,
  1, 3, 3, 1,
  3, 5, 5, 3,
  5, 7, 7, 5,
  1, 3, 3, 1,
  3, 5, 5, 3,
  5, 7, 7, 5 ;

 lat_bnds =
  49.5, 49.5, 50.5, 50.5,
  49.5, 49.5, 50.5, 50.5,
  49.5, 49.5, 50.5, 50.5,
  50.5, 50.5, 51.5, 51.5,
  50.5, 50.5, 51.5, 51.5,
  50.5, 50.5, 51.5, 51.5,
  51.5, 51.5, 52.5, 52.5,
  51.5, 51.5, 52.5, 52.5,
  51.5, 51.5, 52.5, 52.5,
  52.5, 52.5, 53.5, 53.5,
  52.5, 52.5, 53.5, 53.5,
  52.5, 52.5, 53.5, 53.5,
  53.5, 53.5, 54.5, 54.5,
  53.5, 53.5, 54.5, 54.5,
  53.5, 53.5, 54.5, 54.5 ;

 depth =
  1, 106, 11,
  102, 7, 112,
  3, 108, 1.#QNAN,
  104, 9, 114,
  5, 110, 15 ;
}
