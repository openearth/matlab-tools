NetCDF-3 Classic example.nc {

  dimensions:
    lat = 4 ;
    lon = 3 ;
    frtime = UNLIMITED ; (2 currently)
    timelen = 20 ;

  variables:
    // Preference 'PRESERVE_FVD':  false,
    // dimensions consistent with ncBrowse, not with native MATLAB netcdf package.
    single P(frtime,lat,lon), shape = [2 4 3]      :long_name = "pressure at maximum wind" 
      :units = "hectopascals" 
      :valid_range = 0.000000 1500.000000 f
      :_FillValue = -9999.000000 f
    single lat(lat), shape = [4]      :long_name = "latitude" 
      :units = "degrees_north" 
    single lon(lon), shape = [3]      :long_name = "longitude" 
      :units = "degrees_east" 
    int32 frtime(frtime), shape = [2]      :long_name = "forecast time" 
      :units = "hours" 
    char reftime(timelen), shape = [20]      :long_name = "reference time" 
      :units = "text_time" 
    single ScalarVariable([]), shape = [1]
  //global Attributes:
      :history = "created with $Id: netcdf_unidata_only.f90 5822 2012-03-01 14:19:55Z boer_g $ $HeadURL: https://svn.oss.deltares.nl/repos/openearthtools/trunk/fortran/io/netcdf/win32/visual_fortran_6/netcdf_unidata_only.f90 $" 
      :title = "NMC Global Product Set: Pressure at Maximum Wind" 

}
