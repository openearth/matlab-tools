NetCDF-3 Classic d:\checkouts\OpenEarthTools\matlab\io\netcdf\nctools\ncwrite_profile_tutorial_zragged_slow.nc {
dimensions:
	time = 4 ;
	z = 5 ;

variables:
	// Preference 'PRESERVE_FVD':  false,
	// dimensions consistent with ncBrowse, not with native MATLAB netcdf package.
	double time(time), shape = [4]
		time:standard_name = "time" ;
		time:long_name = "time" ;
		time:units = "days since 1970-01-01 00:00:00+00:00" ;
		time:axis = "T" ;
	double z2(time,z), shape = [4 5]
		z2:standard_name = "altitude" ;
		z2:units = "m" ;
		z2:positive = "down" ;
		z2:axis = "Z" ;
		z2:_FillValue = 9.96921e+36 ;
		z2:long_name = "z" ;
		z2:actual_range = 2 18.5 ;
		z2:coordinates = "z2" ;
	double time2(time,z), shape = [4 5]
		time2:standard_name = "time" ;
		time2:long_name = "time" ;
		time2:units = "days since 1970-01-01 00:00:00+00:00" ;
		time2:axis = "T" ;
		time2:coordinates = "z2 time2" ;
	double lon([]), shape = [1]
		lon:standard_name = "longitude" ;
		lon:long_name = "nominal Longitude" ;
		lon:units = "degrees_east" ;
		lon:axis = "X" ;
		lon:_FillValue = 9.96921e+36 ;
		lon:actual_range = 3 3 ;
	double lat([]), shape = [1]
		lat:standard_name = "latitude" ;
		lat:long_name = "nominal Latitude" ;
		lat:units = "degrees_north" ;
		lat:axis = "Y" ;
		lat:_FillValue = 9.96921e+36 ;
		lat:actual_range = 52 52 ;
	double lon1(time), shape = [4]
		lon1:standard_name = "longitude" ;
		lon1:long_name = "drift Longitude" ;
		lon1:units = "degrees_east" ;
		lon1:axis = "X" ;
		lon1:_FillValue = 9.96921e+36 ;
		lon1:actual_range = 2.98287 3.01704 ;
	double lat1(time), shape = [4]
		lat1:standard_name = "latitude" ;
		lat1:long_name = "drift Latitude" ;
		lat1:units = "degrees_north" ;
		lat1:axis = "Y" ;
		lat1:_FillValue = 9.96921e+36 ;
		lat1:actual_range = 51.9911 52.009 ;
	double TSS(time,z), shape = [4 5]
		TSS:standard_name = "mass_concentration_of_suspended_matter_in_sea_water" ;
		TSS:long_name = "TSS" ;
		TSS:units = "kg m-3" ;
		TSS:coordinates = "z2 time2" ;
		TSS:_FillValue = 9.96921e+36 ;
		TSS:actual_range = -1.12559 1.14233 ;
		TSS:xy_comment = "fixed (lat,lon) position, e.g. platform, moored ship" ;
		TSS:z_comment = "varying z levels per profile, e.g. real z positions during of free fall" ;
		TSS:time_comment = "significant time span during one profile, e.g. CTD dangling behind ship for an hour, of slow mechanical lowering" ;

//global attributes:
		:institution = "" ;
		:history = "$HeadURL: https://svn.oss.deltares.nl/repos/openearthtools/trunk/matlab/io/netcdf/nctools/ncwrite_timeseries.m $ $Id: ncwrite_timeseries.m 8921 2013-07-19 06:13:40Z boer_g $" ;
		:featureType = "timeSeriesProfile" ;
		:Conventions = "CF-1.6" ;
		:terms_for_use = "These data can be used freely for research purposes provided that the following source is acknowledged: " ;
		:disclaimer = "This data is made available in the hope that it will be useful, but WITHOUT ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE." ;
		:title = "" ;
		:references = "" ;
		:email = "" ;
		:source = "" ;
		:comment = "" ;
		:version = "" ;
		:time_coverage_start = "20090101T000000" ;
		:time_coverage_end = "20091001T000120" ;
		:geospatial_lat_min = 2.98287 ;
		:geospatial_lat_max = 3.01704 ;
		:geospatial_lon_min = 51.9911 ;
		:geospatial_lon_max = 52.009 ;
		:geospatial_vertical_min = 2 ;
		:geospatial_vertical_max = 18.5 ;


}
