NetCDF-3 Classic nc_cf_grid_write_lat_lon_orthogonal_tutorial.nc {
// The netCDF CF conventions for grids are defined here:
// http://cf-pcmdi.llnl.gov/documents/cf-conventions/1.5/ch05s06.html
// This grid file can be loaded into matlab with nc_cf_grid.m
// To create this netCDF file with Matlab please see nc_cf_grid_write_x_y_orthogonal_tutorial.m

dimensions:
	lon = 3 ;
	lat = 5 ;

variables:
	// Preference 'PRESERVE_FVD':  false,
	// dimensions consistent with ncBrowse, not with native MATLAB netcdf package.
	single lon(lon), shape = [3]
		lon:long_name = "longitude" 
		lon:units = "degrees_east" 
		lon:standard_name = "longitude" 
		lon:actual_range = 2 6 
		lon:grid_mapping = "wgs84" 
	single lat(lat), shape = [5]
		lat:long_name = "latitude" 
		lat:units = "degrees_north" 
		lat:standard_name = "latitude" 
		lat:actual_range = 50 54 
		lat:grid_mapping = "wgs84" 
	int32 wgs84([]), shape = [1]
		wgs84:name = "WGS 84" 
		wgs84:epsg = 4326 
		wgs84:grid_mapping_name = "latitude_longitude" 
		wgs84:semi_major_axis = 6.37814e+006 
		wgs84:semi_minor_axis = 6.35675e+006 
		wgs84:inverse_flattening = 298.257 
		wgs84:comment = "value is equal to EPSG code" 
		wgs84:proj4_params = "+proj=longlat +ellps=WGS84 +datum=WGS84 +no_defs" // non-CF standard required for plotting by ADAGUC
		wgs84:projection_name = "Latitude Longitude"                            // non-CF standard required for plotting by ADAGUC
		wgs84:EPSG_code = "EPSG:4326"                                           // non-CF standard required for plotting by ADAGUC
	single depth(lon,lat), shape = [3 5]
		depth:long_name = "bottom depth" 
		depth:units = "m" 
		depth:_FillValue = NaN f
		depth:actual_range = 1 15 
		depth:coordinates = "lat lon" 
		depth:grid_mapping = "wgs84" 
		depth:standard_name = "sea_floor_depth_below_geoid" 

//global Attributes:
		:title = "" 
		:institution = "" 
		:source = "" 
		:history = "tranformation to netCDF: $HeadURL: https://repos.deltares.nl/repos/OpenEarthTools/trunk/matlab/io/netcdf/nctools/nc_cf_grid_write_lat_lon_orthogonal_tutorial.m $" 
		:references = "" 
		:email = "" 
		:comment = "" 
		:version = "" 
		:Conventions = "CF-1.5" 
		:CF:featureType = "Grid" 
		:terms_for_use = "These data can be used freely for research purposes provided that the following source is acknowledged: " 
		:disclaimer = "This data is made available in the hope that it will be useful, but WITHOUT ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE." 

}
