// Created with Matlab: 2012a 
// with javaclasspath: 
// *  classes 
// *  netcdfAll-4.2.jar 
NetCDF-4 NETCDF4_CLASSIC.nc {

Group / {

  dimensions:
    time = 3 ;
    y = 4 ;
    x = 5 ;

  variables:
    // Preference 'PRESERVE_FVD':  false,
    // dimensions consistent with ncBrowse, not with native MATLAB netcdf package.
    double time(time), shape = [3]
      :units = "seconds since 1970-01-01 00-00-00" 
      :standard_name = "time" 
      :long_name = "time" 
      :_Netcdf4Dimid = 0 d
    double y(y), shape = [4]
      :standard_name = "projection_y_coordinate" 
      :units = "m" 
      :long_name = "y" 
      :_Netcdf4Dimid = 1 d
    double x(x), shape = [5]
      :standard_name = "projection_x_coordinate" 
      :units = "m" 
      :long_name = "x" 
      :_Netcdf4Dimid = 2 d
    single z(time,y,x), shape = [3 4 5]
      :standard_name = "altitude" 
      :units = "m" 
      :long_name = "altitude" 
      :comment = "z = 100*it + 10*iy + ix" 
      :_FillValue = NaN f

  //global Attributes:
      :title = "test file for netCDF format: NETCDF4_CLASSIC" 
      :institution = "Deltares" 
      :source = "Deltares" 
      :history = "$Id: NETCDF_versions_generate.py 7074 2012-07-31 09:31:57Z boer_g $" 
      :references = {''}
      :email = "gerben.deboer@deltares.nl" 
      :comment = {''}
      :version = "Python netCDF4 version 1.0" 
      :Conventions = "CF-1.5" 
      :terms_for_use = "These data can be used freely for research purposes provided that the following source is acknowledged: Deltares" 
      :disclaimer = "This data is made available in the hope that it will be useful, but WITHOUT ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE." 

} End Group /


}
