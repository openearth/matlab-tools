netcdf NETCDF3_64BIT { // format variant: 64bit 
dimensions:
	time = 3 ;
	y = 4 ;
	x = 5 ;
variables:
	double time(time) ;
		time:units = "seconds since 1970-01-01 00-00-00" ;
		time:standard_name = "time" ;
		time:long_name = "time" ;
	double y(y) ;
		y:standard_name = "projection_y_coordinate" ;
		y:units = "m" ;
		y:long_name = "y" ;
	double x(x) ;
		x:standard_name = "projection_x_coordinate" ;
		x:units = "m" ;
		x:long_name = "x" ;
	float z(time, y, x) ;
		z:_FillValue = 1.#QNAN0f ;
		z:standard_name = "altitude" ;
		z:units = "m" ;
		z:long_name = "altitude" ;
		z:comment = "z = 100*it + 10*iy + ix" ;

// global attributes:
		:title = "test file for netCDF format: NETCDF3_64BIT" ;
		:institution = "Deltares" ;
		:source = "Deltares" ;
		:history = "$Id: NETCDF_versions_generate.py 7074 2012-07-31 09:31:57Z boer_g $" ;
		:references = "" ;
		:email = "gerben.deboer@deltares.nl" ;
		:comment = "" ;
		:version = "Python netCDF4 version 1.0" ;
		:Conventions = "CF-1.5" ;
		:terms_for_use = "These data can be used freely for research purposes provided that the following source is acknowledged: Deltares" ;
		:disclaimer = "This data is made available in the hope that it will be useful, but WITHOUT ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE." ;
data:

 time = 0, 1, 2 ;

 y = 0, 1, 2, 3 ;

 x = 0, 1, 2, 3, 4 ;

 z =
  0, 1, 2, 3, 4,
  10, 11, 12, 13, 14,
  20, 21, 22, 23, 24,
  30, 31, 32, 33, 34,
  100, 101, 102, 103, 104,
  110, 111, 112, 113, 114,
  120, 121, 122, 123, 124,
  130, 131, 132, 133, 134,
  200, 201, 202, 203, 204,
  210, 211, 212, 213, 214,
  220, 221, 222, 223, 224,
  230, 231, 232, 233, 234 ;
}
