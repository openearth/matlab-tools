// The netCDF CF conventions for grids are defined here:
// http://cf-pcmdi.llnl.gov/documents/cf-conventions/1.6/ch05s06.html
// This grid file can be loaded into matlab with nc_cf_grid.m and d3d_qp.m
// To create this netCDF file with Matlab please see nc_cf_grid_write_x_y_orthogonal_tutorial
NetCDF-3 Classic nc_cf_grid_write_x_y_orthogonal_tutorial.nc {

  dimensions:
    x = 3 ;
    y = 5 ;
    time = 1 ;

  variables:
    // Preference 'PRESERVE_FVD':  false,
    // dimensions consistent with ncBrowse, not with native MATLAB netcdf package.
    single x(x), shape = [3]
      :long_name = "x Rijksdriehoek" 
      :units = "m" 
      :standard_name = "projection_x_coordinate" 
      :actual_range = 400000 600000 
      :grid_mapping = "epsg" 
    single y(y), shape = [5]
      :long_name = "y Rijksdriehoek" 
      :units = "m" 
      :standard_name = "projection_y_coordinate" 
      :actual_range = 5.5e+06 5.9e+06 
      :grid_mapping = "epsg" 
    int32 epsg([]), shape = [1]
      :name = "WGS 84 / UTM zone 31N" 
      :epsg = 32631 
      :epsg_name = "Transverse Mercator" 
      :grid_mapping_name = "transverse_mercator" 
      :semi_major_axis = 6.37814e+06 
      :semi_minor_axis = 6.35675e+06 
      :inverse_flattening = 298.257 
      :latitude_of_projection_origin = 0 
      :longitude_of_projection_origin = 3 
      :false_easting = 500000 
      :false_northing = 0 
      :scale_factor_at_projection_origin = 0.9996 
      :proj4_params = "+proj=utm +zone=31 +ellps=WGS84 +datum=WGS84 +units=m +no_defs " 
      :EPSG_code = "EPSG:32631" 
      :projection_name = "WGS 84 / UTM zone 31N" 
      :wkt = "" 
      :comment = "value is equal to EPSG code" 
    single lon(x,y), shape = [3 5]
      :long_name = "longitude" 
      :units = "degrees_east" 
      :standard_name = "longitude" 
      :actual_range = 1.50155 4.49845 
      :coordinates = "lat lon" 
      :grid_mapping = "wgs84" 
    single lat(x,y), shape = [3 5]
      :long_name = "latitude" 
      :units = "degrees_north" 
      :standard_name = "latitude" 
      :actual_range = 49.6443 53.2493 
      :coordinates = "lat lon" 
      :grid_mapping = "wgs84" 
    int32 wgs84([]), shape = [1]
      :name = "WGS 84" 
      :epsg = 4326 
      :grid_mapping_name = "latitude_longitude" 
      :semi_major_axis = 6.37814e+06 
      :semi_minor_axis = 6.35675e+06 
      :inverse_flattening = 298.257 
      :proj4_params = "+proj=longlat +ellps=WGS84 +datum=WGS84 +no_defs " 
      :EPSG_code = "EPSG:4326" 
      :projection_name = "Latitude Longitude" 
      :wkt = "" 
      :comment = "value is equal to EPSG code" 
    double time(time), shape = [1]
      :long_name = "time" 
      :units = "days since 1970-01-01 00:00:00 +00:00" 
      :standard_name = "time" 
      :actual_range = 15833.7 15833.7 
    single depth(time,x,y), shape = [1 3 5]
      :long_name = "bottom depth" 
      :units = "m" 
      :_FillValue = NaN f
      :actual_range = 1 114 
      :coordinates = "lat lon" 
      :grid_mapping = "epsg" 
      :standard_name = "sea_floor_depth_below_geoid" 

  //global Attributes:
      :title = "" 
      :institution = "" 
      :source = "" 
      :history = "tranformation to netCDF: $HeadURL: https://svn.oss.deltares.nl/repos/openearthtools/trunk/matlab/io/netcdf/nctools/nc_cf_grid_write_x_y_orthogonal_tutorial.m $" 
      :references = "" 
      :email = "" 
      :comment = "" 
      :version = "" 
      :Conventions = "CF-1.5" 
      :CF:featureType = "Grid" 
      :terms_for_use = "These data can be used freely for research purposes provided that the following source is acknowledged: " 
      :disclaimer = "This data is made available in the hope that it will be useful, but WITHOUT ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE." 


}
