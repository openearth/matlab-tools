NetCDF-3 Classic nc_cf_grid_write_lat_lon_orthogonal_tutorial.nc {

  dimensions:
    lon = 3 ;
    lat = 5 ;
    vertices = 2 ;
    time = 1 ;

  variables:
    // Preference 'PRESERVE_FVD':  false,
    // dimensions consistent with ncBrowse, not with native MATLAB netcdf package.
    double time(time), shape = [1]
      :standard_name = "time" 
      :long_name = "time" 
      :units = "days since 1970-01-01 00:00:00 +00:00" 
      :actual_range = 15833.7 15833.7 
    single lon(lon), shape = [3]
      :long_name = "longitude" 
      :units = "degrees_east" 
      :standard_name = "longitude" 
      :actual_range = 2 6 
      :grid_mapping = "wgs84" 
      :bounds = "lonbounds" 
    single lonbounds(lon,vertices), shape = [3 2]
      :long_name = "longitude vertices" 
      :units = "degrees_east" 
      :standard_name = "longitude" 
      :actual_range = 1 7 
      :grid_mapping = "wgs84" 
    single lat(lat), shape = [5]
      :long_name = "latitude" 
      :units = "degrees_north" 
      :standard_name = "latitude" 
      :actual_range = 50 54 
      :grid_mapping = "wgs84" 
      :bounds = "latbounds" 
    single latbounds(lat,vertices), shape = [5 2]
      :long_name = "latitude vertices" 
      :units = "degrees_north" 
      :standard_name = "latitude" 
      :actual_range = 49.5 54.5 
      :grid_mapping = "wgs84" 
    int32 wgs84([]), shape = [1]
      :name = "WGS 84" 
      :epsg = 4326 
      :grid_mapping_name = "latitude_longitude" 
      :semi_major_axis = 6.37814e+06 
      :semi_minor_axis = 6.35675e+06 
      :inverse_flattening = 298.257 
      :comment = "value is equal to EPSG code" 
      :proj4_params = "+proj=longlat +ellps=WGS84 +datum=WGS84 +no_defs" 
      :projection_name = "Latitude Longitude" 
      :EPSG_code = "EPSG:4326" 
    single depth(time,lon,lat), shape = [1 3 5]
      :long_name = "bottom depth" 
      :units = "m" 
      :_FillValue = NaN f
      :actual_range = 1 114 
      :coordinates = "lat lon" 
      :grid_mapping = "wgs84" 
      :standard_name = "sea_floor_depth_below_geoid" 

  //global Attributes:
      :title = "" 
      :institution = "" 
      :source = "" 
      :history = "tranformation to netCDF: $HeadURL: https://svn.oss.deltares.nl/repos/openearthtools/trunk/matlab/io/netcdf/nctools/nc_cf_grid_write_lat_lon_orthogonal_tutorial.m $" 
      :references = "" 
      :email = "" 
      :comment = "" 
      :version = "" 
      :Conventions = "CF-1.5" 
      :CF:featureType = "Grid" 
      :terms_for_use = "These data can be used freely for research purposes provided that the following source is acknowledged: " 
      :disclaimer = "This data is made available in the hope that it will be useful, but WITHOUT ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE." 


}
