NetCDF-3 Classic ncwritetutorial_grid_lat_lon_curvilinear.nc {

  dimensions:
    col = 3 ;
    row = 5 ;
    time = 1 ;
    bounds = 4 ;

  variables:
    // Preference 'PRESERVE_FVD':  false,
    // dimensions consistent with ncBrowse, not with native MATLAB netcdf package.
    double time(time), shape = [1]
      :standard_name = "time" 
      :long_name = "time" 
      :units = "days since 1970-01-01 00:00:00+08:00" 
      :axis = "T" 
    double longitude(row,col), shape = [5 3]
      :standard_name = "longitude" 
      :long_name = "Longitude" 
      :units = "degrees_east" 
      :axis = "X" 
      :_FillValue = NaN 
      :coordinates = "longitude latitude" 
      :actual_range = 2.78657 8.94889 
      :bounds = "longitude_bounds" 
    double latitude(row,col), shape = [5 3]
      :standard_name = "latitude" 
      :long_name = "Latitude" 
      :units = "degrees_north" 
      :axis = "Y" 
      :_FillValue = NaN 
      :coordinates = "longitude latitude" 
      :actual_range = 48.8618 55.8107 
      :bounds = "latitude_bounds" 
    double longitude_bounds(row,col,bounds), shape = [5 3 4]
      :standard_name = "longitude" 
      :long_name = "Longitude" 
      :units = "degrees_east" 
      :axis = "X" 
      :_FillValue = NaN 
      :actual_range = 2.78657 8.94889 
    double latitude_bounds(row,col,bounds), shape = [5 3 4]
      :standard_name = "latitude" 
      :long_name = "Latitude" 
      :units = "degrees_north" 
      :axis = "Y" 
      :_FillValue = NaN 
      :actual_range = 48.8618 55.8107 
    double depth(time,row,col), shape = [1 5 3]
      :standard_name = "sea_floor_depth_below_geoid" 
      :long_name = "bottom depth" 
      :units = "m" 
      :_FillValue = NaN 
      :coordinates = "longitude latitude" 
      :actual_range = 1 114 

  //global Attributes:
      :title = "" 
      :institution = "Deltares" 
      :source = "" 
      :history = "$HeadURL: https://svn.oss.deltares.nl/repos/openearthtools/trunk/matlab/io/netcdf/nctools/ncwritetutorial_grid_lat_lon_curvilinear.m $ $Id: ncwritetutorial_grid.m 8596 2013-05-08 16:08:39Z boer_g $" 
      :references = "http://svn.oss.deltares.nl" 
      :email = "" 
      :featureType = "grid" 
      :comment = "" 
      :version = "" 
      :Conventions = "CF-1.6" 
      :terms_for_use = "These data can be used freely for research purposes provided that the following source is acknowledged: Deltares" 
      :disclaimer = "This data is made available in the hope that it will be useful, but WITHOUT ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE." 


}
