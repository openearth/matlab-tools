netcdf netCDF4_tutorial_grid_lat_lon_orthogonal {
dimensions:
	lat = 5 ;
	lon = 3 ;
	time = 1 ;
	bounds = 2 ;
variables:
	double time(time) ;
		time:standard_name = "time" ;
		time:long_name = "time" ;
		time:units = "seconds since 1970-01-01 00-00-00" ;
		time:axis = "T" ;
	double lat(lat) ;
		lat:_FillValue = NaN ;
		lat:standard_name = "latitude" ;
		lat:long_name = "Latitude" ;
		lat:units = "degrees_north" ;
		lat:axis = "Y" ;
		lat:grid_mapping = "projection" ;
		lat:actual_range = 50., 54. ;
		lat:bounds = "lat_bnds" ;
	double lon(lon) ;
		lon:_FillValue = NaN ;
		lon:standard_name = "longitude" ;
		lon:long_name = "Longitude" ;
		lon:units = "degrees_east" ;
		lon:axis = "X" ;
		lon:grid_mapping = "projection" ;
		lon:actual_range = 1.5, 3.5 ;
		lon:bounds = "lon_bnds" ;
	int projection ;
		projection:name = "WGS 84" ;
		projection:epsg = 4326. ;
		projection:grid_mapping_name = "latitude_longitude" ;
		projection:semi_major_axis = 6378137. ;
		projection:semi_minor_axis = 6356752.31424783 ;
		projection:inverse_flattening = 298.2572236 ;
		projection:proj4_params = "+proj=longlat +ellps=WGS84 +datum=WGS84 +no_defs" ;
		projection:projection_name = "Latitude Longitude" ;
		projection:EPSG_code = "EPSG:4326" ;
	double lon_bnds(bounds, lon) ;
		lon_bnds:_FillValue = NaN ;
		lon_bnds:standard_name = "longitude" ;
		lon_bnds:long_name = "Longitude bounds" ;
		lon_bnds:units = "degrees_east" ;
		lon_bnds:actual_range = 1., 4. ;
	double lat_bnds(bounds, lat) ;
		lat_bnds:_FillValue = NaN ;
		lat_bnds:standard_name = "latitude" ;
		lat_bnds:long_name = "Latitude bounds" ;
		lat_bnds:units = "degrees_north" ;
		lat_bnds:actual_range = 49.5, 54.5 ;
	float depth(time, lat, lon) ;
		depth:_FillValue = NaNf ;
		depth:standard_name = "sea_floor_depth_below_geoid" ;
		depth:long_name = "bottom depth" ;
		depth:units = "m" ;
		depth:positive = "up" ;
		depth:actual_range = 1., 114. ;
		depth:grid_mapping = "projection" ;
		depth:coordinates = "lat lon" ;

// global attributes:
		:title = "ncwritetutorial_grid_lat_lon_orthogonal" ;
		:institution = "Deltares" ;
		:source = "" ;
		:history = "$HeadURL: https://svn.oss.deltares.nl/repos/openearthtools/trunk/matlab/io/netcdf/nctools/ncwritetutorial_grid_lat_lon_curvilinear.m $ $Id: ncwritetutorial_grid_lat_lon_curvilinear.m 8901 2013-07-09 06:51:31Z boer_g $" ;
		:references = "http://svn.oss.deltares.nl" ;
		:email = "" ;
		:featureType = "Grid" ;
		:comment = "" ;
		:version = "beta" ;
		:Conventions = "CF-1.6" ;
		:terms_for_use = "These data can be used freely for research purposes provided that the following source is acknowledged: Deltares" ;
		:disclaimer = "This data is made available in the hope that it will be useful, but WITHOUT ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE." ;
data:

 time = 946681200 ;

 lat = 50, 51, 52, 53, 54 ;

 lon = 1.5, 2.5, 3.5 ;

 projection = _ ;

 lon_bnds =
  1, 2, 2,
  3, 3, 4 ;

 lat_bnds =
  49.5, 50.5, 50.5, 51.5, 51.5,
  52.5, 52.5, 53.5, 53.5, 54.5 ;

 depth =
  1, 106, 11,
  102, 7, 112,
  3, 108, _,
  104, 9, 114,
  5, 110, 15 ;
}
