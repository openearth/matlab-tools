NetCDF-3 Classic d:\checkouts\OpenEarthTools\matlab\io\netcdf\nctools\ncwritetutorial_trajectory.nc {
dimensions:
	time = 365 ;

variables:
	// Preference 'PRESERVE_FVD':  false,
	// dimensions consistent with ncBrowse, not with native MATLAB netcdf package.
	double time(time), shape = [365]
		time:standard_name = "time" ;
		time:long_name = "time" ;
		time:units = "days since 1970-01-01 00:00:00+00:00" ;
		time:axis = "T" ;
	double lon(time), shape = [365]
		lon:standard_name = "longitude" ;
		lon:long_name = "Longitude" ;
		lon:units = "degrees_east" ;
		lon:axis = "X" ;
		lon:_FillValue = 9.96921e+36 ;
		lon:actual_range = 1.00007 5 ;
	double lat(time), shape = [365]
		lat:standard_name = "latitude" ;
		lat:long_name = "Latitude" ;
		lat:units = "degrees_north" ;
		lat:axis = "Y" ;
		lat:_FillValue = 9.96921e+36 ;
		lat:actual_range = 51 53 ;
	double z(time), shape = [365]
		z:standard_name = "altitude" ;
		z:long_name = "z" ;
		z:units = "m" ;
		z:positive = "down" ;
		z:axis = "Z" ;
		z:_FillValue = 9.96921e+36 ;
		z:actual_range = -0.999963 1 ;
	double TSS(time), shape = [365]
		TSS:standard_name = "mass_concentration_of_suspended_matter_in_sea_water" ;
		TSS:long_name = "TSS" ;
		TSS:units = "kg m-3" ;
		TSS:coordinates = "lat lon" ;
		TSS:_FillValue = 9.96921e+36 ;
		TSS:actual_range = 1 4.99993 ;

//global attributes:
		:title = "" ;
		:institution = "" ;
		:source = "" ;
		:history = "$HeadURL: https://svn.oss.deltares.nl/repos/openearthtools/trunk/matlab/io/netcdf/nctools/ncwritetutorial_timeseries.m $ $Id: ncwritetutorial_timeseries.m 8921 2013-07-19 06:13:40Z boer_g $" ;
		:references = "" ;
		:email = "" ;
		:featureType = "timeSeries" ;
		:comment = "" ;
		:version = "" ;
		:Conventions = "CF-1.6" ;
		:terms_for_use = "These data can be used freely for research purposes provided that the following source is acknowledged: " ;
		:disclaimer = "This data is made available in the hope that it will be useful, but WITHOUT ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE." ;


}
