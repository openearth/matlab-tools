// The netCDF-CF conventions for grids are defined here:
// http://cf-pcmdi.llnl.gov/documents/cf-conventions/
// This grid file can be loaded into matlab with QuickPlot (d3d_qp.m) and ADAGUC.knmi.nl.
// To create this netCDF file with Matlab please see ncwritetutorial_grid_x_y_curvilinear
NetCDF-3 Classic ncwritetutorial_grid_x_y_curvilinear.nc {

  dimensions:
    col = 3 ;
    row = 5 ;
    time = 1 ;
    bounds = 4 ;

  variables:
    // Preference 'PRESERVE_FVD':  false,
    // dimensions consistent with ncBrowse, not with native MATLAB netcdf package.
    double time(time), shape = [1]
      :standard_name = "time" 
      :long_name = "time" 
      :units = "days since 1970-01-01 00:00:00+08:00" 
      :axis = "T" 
    double x(row,col), shape = [5 3]
      :standard_name = "projection_x_coordinate" 
      :long_name = "Easting" 
      :units = "m" 
      :axis = "X" 
      :_FillValue = NaN 
      :grid_mapping = "epsg" 
      :actual_range = 314268 853681 
      :bounds = "lon_bnds" 
    double y(row,col), shape = [5 3]
      :standard_name = "projection_y_coordinate" 
      :long_name = "Northing" 
      :units = "m" 
      :axis = "Y" 
      :_FillValue = NaN 
      :grid_mapping = "epsg" 
      :actual_range = 5.39144e+06 6.13469e+06 
      :bounds = "lat_bnds" 
    double lon(row,col), shape = [5 3]
      :standard_name = "longitude" 
      :long_name = "Longitude" 
      :units = "degrees_east" 
      :axis = "X" 
      :_FillValue = NaN 
      :grid_mapping = "wgs84" 
      :actual_range = 0.125 7.875 
      :bounds = "lon_bnds" 
    double lat(row,col), shape = [5 3]
      :standard_name = "latitude" 
      :long_name = "Latitude" 
      :units = "degrees_north" 
      :axis = "Y" 
      :_FillValue = NaN 
      :grid_mapping = "wgs84" 
      :actual_range = 48.65 55.35 
      :bounds = "lat_bnds" 
    int32 epsg([]), shape = [1]
      :name = "WGS 84 / UTM zone 31N" 
      :epsg = 32631 
      :epsg_name = "Transverse Mercator" 
      :grid_mapping_name = "transverse_mercator" 
      :semi_major_axis = 6.37814e+06 
      :semi_minor_axis = 6.35675e+06 
      :inverse_flattening = 298.257 
      :latitude_of_projection_origin = 0 
      :longitude_of_projection_origin = 3 
      :false_easting = 500000 
      :false_northing = 0 
      :scale_factor_at_projection_origin = 0.9996 
      :proj4_params = "+proj=utm +zone=31 +ellps=WGS84 +datum=WGS84 +units=m +no_defs " 
      :EPSG_code = "EPSG:32631" 
      :projection_name = "WGS 84 / UTM zone 31N" 
      :wkt = "" 
      :comment = "value is equal to EPSG code" 
    int32 wgs84([]), shape = [1]
      :name = "WGS 84" 
      :epsg = 4326 
      :grid_mapping_name = "latitude_longitude" 
      :semi_major_axis = 6.37814e+06 
      :semi_minor_axis = 6.35675e+06 
      :inverse_flattening = 298.257 
      :proj4_params = "+proj=longlat +ellps=WGS84 +datum=WGS84 +no_defs" 
      :EPSG_code = "EPSG:4326" 
      :projection_name = "Latitude Longitude" 
      :wkt = "" 
      :comment = "value is equal to EPSG code" 
    double x_bnds(row,col,bounds), shape = [5 3 4]
      :standard_name = "projection_x_coordinate" 
      :long_name = "Easting bounds" 
      :units = "m" 
      :_FillValue = NaN 
      :actual_range = 111663 1.07896e+06 
    double y_bnds(row,col,bounds), shape = [5 3 4]
      :standard_name = "projection_y_coordinate" 
      :long_name = "Northing bounds" 
      :units = "m" 
      :_FillValue = NaN 
      :actual_range = 5.26121e+06 6.26352e+06 
    double lon_bnds(row,col,bounds), shape = [5 3 4]
      :standard_name = "longitude" 
      :long_name = "Longitude bounds" 
      :units = "degrees_east" 
      :_FillValue = NaN 
      :actual_range = -3 11 
    double lat_bnds(row,col,bounds), shape = [5 3 4]
      :standard_name = "latitude" 
      :long_name = "Latitude bounds" 
      :units = "degrees_north" 
      :_FillValue = NaN 
      :actual_range = 47.5 56.5 
    double depth(time,row,col), shape = [1 5 3]
      :standard_name = "sea_floor_depth_below_geoid" 
      :long_name = "bottom depth" 
      :units = "m" 
      :_FillValue = NaN 
      :actual_range = 1 114 
      :grid_mapping = "epsg" 
      :coordinates = "lat lon" 

  //global Attributes:
      :title = "ncwritetutorial_grid_x_y_curvilinear" 
      :institution = "Deltares" 
      :source = "" 
      :history = "$HeadURL: https://svn.oss.deltares.nl/repos/openearthtools/trunk/matlab/io/netcdf/nctools/ncwritetutorial_grid_x_y_curvilinear.m $ $Id: ncwritetutorial_grid_x_y_curvilinear.m 8831 2013-06-19 08:05:18Z boer_g $" 
      :references = "http://svn.oss.deltares.nl" 
      :email = "" 
      :featureType = "grid" 
      :comment = "" 
      :version = "" 
      :Conventions = "CF-1.6" 
      :terms_for_use = "These data can be used freely for research purposes provided that the following source is acknowledged: Deltares" 
      :disclaimer = "This data is made available in the hope that it will be useful, but WITHOUT ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE." 
      :time_coverage_start = "2000-01-01T00:00" 
      :time_coverage_end = "2000-01-01T00:00" 


}
