// The netCDF CF conventions for grids are defined here:
// http://cf-pcmdi.llnl.gov/documents/cf-conventions/1.6/ch05s06.html
// This grid file can be loaded into matlab with nc_cf_grid.m and d3d_qp.m
// To create this netCDF file with Matlab please see nc_cf_grid_write_lat_lon_curvilinear_tutorial
NetCDF-3 Classic nc_cf_grid_write_lat_lon_curvilinear_tutorial.nc {

  dimensions:
    col = 3 ;
    row = 5 ;
    vertices = 4 ;
    time = 1 ;

  variables:
    // Preference 'PRESERVE_FVD':  false,
    // dimensions consistent with ncBrowse, not with native MATLAB netcdf package.
    single lon(col,row), shape = [3 5]
      :long_name = "longitude" 
      :units = "degrees_east" 
      :standard_name = "longitude" 
      :actual_range = 2.78657 8.94889 
      :coordinates = "lat lon" 
      :grid_mapping = "wgs84" 
      :bounds = "lonbounds" 
    single lonbounds(col,row,vertices), shape = [3 5 4]
      :long_name = "longitude vertices" 
      :units = "degrees_east" 
      :standard_name = "longitude" 
      :actual_range = 1.35355 10.5 
      :coordinates = "lat lon" 
      :grid_mapping = "wgs84" 
    single lat(col,row), shape = [3 5]
      :long_name = "latitude" 
      :units = "degrees_north" 
      :standard_name = "latitude" 
      :actual_range = 48.8618 55.8107 
      :coordinates = "lat lon" 
      :grid_mapping = "wgs84" 
      :bounds = "latbounds" 
    single latbounds(col,row,vertices), shape = [3 5 4]
      :long_name = "latitude vertices" 
      :units = "degrees_north" 
      :standard_name = "latitude" 
      :actual_range = 47.75 56.9749 
      :coordinates = "lat lon" 
      :grid_mapping = "wgs84" 
    int32 wgs84([]), shape = [1]
      :name = "WGS 84" 
      :epsg = 4326 
      :grid_mapping_name = "latitude_longitude" 
      :semi_major_axis = 6.37814e+06 
      :semi_minor_axis = 6.35675e+06 
      :inverse_flattening = 298.257 
      :comment = "value is equal to EPSG code" 
      :proj4_params = "+proj=longlat +ellps=WGS84 +datum=WGS84 +no_defs" 
      :projection_name = "Latitude Longitude" 
      :EPSG_code = "EPSG:4326" 
    double time(time), shape = [1]
      :long_name = "time" 
      :units = "days since 1970-01-01 00:00:00 +00:00" 
      :standard_name = "time" 
      :actual_range = 15833.7 15833.7 
    single depth(time,col,row), shape = [1 3 5]
      :long_name = "bottom depth" 
      :units = "m" 
      :_FillValue = NaN f
      :actual_range = 1 114 
      :coordinates = "lat lon" 
      :grid_mapping = "wgs84" 
      :standard_name = "sea_floor_depth_below_geoid" 

  //global Attributes:
      :title = "" 
      :institution = "" 
      :source = "" 
      :history = "tranformation to netCDF: $HeadURL: https://svn.oss.deltares.nl/repos/openearthtools/trunk/matlab/io/netcdf/nctools/nc_cf_grid_write_lat_lon_curvilinear_tutorial.m $" 
      :references = "" 
      :email = "" 
      :comment = "" 
      :version = "" 
      :Conventions = "CF-1.5" 
      :CF:featureType = "Grid" 
      :terms_for_use = "These data can be used freely for research purposes provided that the following source is acknowledged: " 
      :disclaimer = "This data is made available in the hope that it will be useful, but WITHOUT ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE." 


}
