// The netCDF-CF conventions for grids are defined here:
// http://cf-pcmdi.llnl.gov/documents/cf-conventions/
// This grid file can be loaded into matlab with QuickPlot (d3d_qp.m) and ADAGUC.knmi.nl.
// To create this netCDF file with Matlab please see nc_cf_grid_write_lat_lon_orthogonal_tutorial
NetCDF-3 Classic nc_cf_grid_write_lat_lon_orthogonal_tutorial.nc {

  dimensions:
    lon = 3 ;
    lat = 5 ;
    time = 1 ;
    bounds = 2 ;

  variables:
    // Preference 'PRESERVE_FVD':  false,
    // dimensions consistent with ncBrowse, not with native MATLAB netcdf package.
    double time(time), shape = [1]
      :standard_name = "time" 
      :long_name = "time" 
      :units = "days since 1970-01-01 00:00:00 +08:00" 
      :axis = "T" 
    double lon(lon), shape = [3]
      :standard_name = "longitude" 
      :long_name = "Longitude" 
      :units = "degrees_east" 
      :axis = "X" 
      :grid_mapping = "wgs84" 
      :actual_range = 2 6 
      :bounds = "lon_bnds" 
    double lat(lat), shape = [5]
      :standard_name = "latitude" 
      :long_name = "Latitude" 
      :units = "degrees_north" 
      :axis = "Y" 
      :grid_mapping = "wgs84" 
      :actual_range = 50 54 
      :bounds = "lat_bnds" 
    int32 wgs84([]), shape = [1]
      :name = "WGS 84" 
      :epsg = 4326 
      :grid_mapping_name = "latitude_longitude" 
      :semi_major_axis = 6.37814e+06 
      :semi_minor_axis = 6.35675e+06 
      :inverse_flattening = 298.257 
      :comment = "value is equal to EPSG code" 
      :proj4_params = "+proj=longlat +ellps=WGS84 +datum=WGS84 +no_defs" 
      :projection_name = "Latitude Longitude" 
      :EPSG_code = "EPSG:4326" 
    double lon_bnds(lon,bounds), shape = [3 2]
      :standard_name = "longitude" 
      :long_name = "Longitude bounds" 
      :units = "degrees_east" 
      :actual_range = 1 7 
    double lat_bnds(lat,bounds), shape = [5 2]
      :standard_name = "latitude" 
      :long_name = "Latitude bounds" 
      :units = "degrees_north" 
      :actual_range = 49.5 54.5 
    double depth(time,lat,lon), shape = [1 5 3]
      :standard_name = "sea_floor_depth_below_geoid" 
      :long_name = "bottom depth" 
      :units = "m" 
      :actual_range = 1 114 
      :grid_mapping = "wgs84" 

  //global Attributes:
      :title = "nc_cf_grid_write_lat_lon_orthogonal_tutorial" 
      :institution = "Deltares" 
      :source = "" 
      :history = "$HeadURL: https://svn.oss.deltares.nl/repos/openearthtools/trunk/matlab/io/netcdf/nctools/nc_cf_grid_write_lat_lon_orthogonal_tutorial.m $ $Id: nc_cf_grid_write_lat_lon_orthogonal_tutorial.m 8825 2013-06-18 14:19:32Z boer_g $" 
      :references = "http://svn.oss.deltares.nl" 
      :email = "" 
      :featureType = "grid" 
      :comment = "" 
      :version = "" 
      :Conventions = "CF-1.6" 
      :terms_for_use = "These data can be used freely for research purposes provided that the following source is acknowledged: Deltares" 
      :disclaimer = "This data is made available in the hope that it will be useful, but WITHOUT ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE." 
      :time_coverage_start = "2013-06-18T21:55" 
      :time_coverage_end = "2013-06-18T21:55" 


}
