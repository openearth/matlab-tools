NetCDF F:\checkouts\OpenEarthTools\matlab\io\netcdf\nctools\nc_cf_grid_write_x_y_curvilinear_tutorial.nc {

// The netCDF CF conventions for grids are defined here:
// http://cf-pcmdi.llnl.gov/documents/cf-conventions/1.5/ch05s06.html
// This grid file can be loaded into matlab with nc_cf_grid.m
// To create this netCDF file with Matlab please see nc_cf_grid_write_x_y_curvilinear_tutorial.m

dimensions:
	col = 3 ;
	row = 5 ;

variables:
	// Preference 'PRESERVE_FVD':  false,
	// dimensions consistent with ncBrowse, not with native MATLAB netcdf package.
	single x(col,row), shape = [3 5]
		x:long_name = "x Rijksdriehoek" 
		x:units = "m" 
		x:standard_name = "projection_x_coordinate" 
		x:actual_range = 481128 929333 
		x:coordinates = "lat lon" 
		x:grid_mapping = "epsg" 
	single y(col,row), shape = [3 5]
		y:long_name = "y Rijksdriehoek" 
		y:units = "m" 
		y:standard_name = "projection_y_coordinate" 
		y:actual_range = 5.46907e+006 6.2314e+006 
		y:coordinates = "lat lon" 
		y:grid_mapping = "epsg" 
	int32 epsg([]), shape = [1]
		epsg:name = "WGS 84 / UTM zone 31N" 
		epsg:epsg = 32631 
		epsg:epsg_name = "Transverse Mercator" 
		epsg:grid_mapping_name = "transverse_mercator" 
		epsg:semi_major_axis = 6.37814e+006 
		epsg:semi_minor_axis = 6.35675e+006 
		epsg:inverse_flattening = 298.257 
		epsg:latitude_of_projection_origin = 0 
		epsg:longitude_of_projection_origin = 3 
		epsg:false_easting = 500000 
		epsg:false_northing = 0 
		epsg:scale_factor_at_projection_origin = 0.9996 
		epsg:proj4_params = "+proj=utm +zone=31 +ellps=WGS84 +datum=WGS84 +units=m +no_defs " 
		epsg:EPSG_code = "EPSG:32631" 
		epsg:projection_name = "WGS 84 / UTM zone 31N" 
		epsg:wkt = "PROJCS["WGS 84 / UTM zone 31N",
    GEOGCS["WGS 84",
        DATUM["WGS_1984",
            SPHEROID["WGS 84",6378137,298.257223563,
                AUTHORITY["EPSG","7030"]],
            AUTHORITY["EPSG","6326"]],
        PRIMEM["Greenwich",0,
            AUTHORITY["EPSG","8901"]],
        UNIT["degree",0.01745329251994328,
            AUTHORITY["EPSG","9122"]],
        AUTHORITY["EPSG","4326"]],
    UNIT["metre",1,
        AUTHORITY["EPSG","9001"]],
    PROJECTION["Transverse_Mercator"],
    PARAMETER["latitude_of_origin",0],
    PARAMETER["central_meridian",3],
    PARAMETER["scale_factor",0.9996],
    PARAMETER["false_easting",500000],
    PARAMETER["false_northing",0],
    AUTHORITY["EPSG","32631"],
    AXIS["Easting",EAST],
    AXIS["Northing",NORTH]]" 
		epsg:comment = "value is equal to EPSG code" 
	single lon(col,row), shape = [3 5]
		lon:long_name = "longitude" 
		lon:units = "degrees_east" 
		lon:standard_name = "longitude" 
		lon:actual_range = 2.70711 9 
		lon:coordinates = "x y" 
		lon:grid_mapping = "wgs84" 
	single lat(col,row), shape = [3 5]
		lat:long_name = "latitude" 
		lat:units = "degrees_north" 
		lat:standard_name = "latitude" 
		lat:actual_range = 49.2235 56.1213 
		lat:coordinates = "x y" 
		lat:grid_mapping = "wgs84" 
	int32 wgs84([]), shape = [1]
		wgs84:name = "WGS 84" 
		wgs84:epsg = 4326 
		wgs84:grid_mapping_name = "latitude_longitude" 
		wgs84:semi_major_axis = 6.37814e+006 
		wgs84:semi_minor_axis = 6.35675e+006 
		wgs84:inverse_flattening = 298.257 
		wgs84:proj4_params = "+proj=longlat +ellps=WGS84 +datum=WGS84 +no_defs " 
		wgs84:EPSG_code = "EPSG:4326" 
		wgs84:projection_name = "Latitude Longitude" 
		wgs84:wkt = "GEOGCS["WGS 84",
    DATUM["WGS_1984",
        SPHEROID["WGS 84",6378137,298.257223563,
            AUTHORITY["EPSG","7030"]],
        AUTHORITY["EPSG","6326"]],
    PRIMEM["Greenwich",0,
        AUTHORITY["EPSG","8901"]],
    UNIT["degree",0.01745329251994328,
        AUTHORITY["EPSG","9122"]],
    AUTHORITY["EPSG","4326"]]" 
		wgs84:comment = "value is equal to EPSG code" 
	single depth(col,row), shape = [3 5]
		depth:long_name = "bottom depth" 
		depth:units = "m" 
		depth:_FillValue = NaN f
		depth:actual_range = 1 15 
		depth:coordinates = "lat lon" 
		depth:coordinates2 = "x y" 
		depth:grid_mapping = "wgs84" 
		depth:standard_name = "sea_floor_depth_below_geoid" 

//global Attributes:
		:title = " " 
		:institution = " " 
		:source = " " 
		:history = "tranformation to netCDF: $HeadURL: https://repos.deltares.nl/repos/OpenEarthTools/trunk/matlab/io/netcdf/nctools/nc_cf_grid_write_x_y_curvilinear_tutorial.m $" 
		:references = " " 
		:email = " " 
		:comment = " " 
		:version = " " 
		:Conventions = "CF-1.5" 
		:CF:featureType = "Grid" 
		:terms_for_use = "These data can be used freely for research purposes provided that the following source is acknowledged: " 
		:disclaimer = "This data is made available in the hope that it will be useful, but WITHOUT ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE." 

}
